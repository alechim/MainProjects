Make;Model;MPG;Cylinders;Displacement;Horsepower;Weight;Year;Origin
Ford;Mustang;25.5;6;3000;350;3000;2022;USA
Chevrolet;Camaro;24.8;8;3500;400;3200;2023;USA
Toyota;Corolla;35.2;4;2000;150;2500;2023;Japan
Honda;Accord;31.5;6;2800;300;2900;2022;Japan
BMW;M3;27.8;6;3200;380;3300;2022;Germany
Mercedes-Benz;C-Class;29.6;4;2500;280;2800;2023;Germany
Hyundai;Elantra;33.1;4;2200;160;2700;2023;South Korea
Nissan;Altima;30.2;6;2900;270;3000;2022;Japan
Audi;A4;28.7;4;2700;300;2900;2022;Germany
Lexus;ES;32.5;6;3100;320;3200;2023;Japan
Kia;Optima;29.8;4;2600;180;2800;2022;South Korea
Subaru;Legacy;30.9;6;3000;250;2900;2023;Japan
Volkswagen;Passat;31.8;4;2800;220;3000;2022;Germany
Mazda;6;28.5;4;2700;200;2800;2022;Japan
Tesla;Model 3;140.5;0;0;450;3500;2023;USA
Ford;Focus;30.0;4;2200;160;2700;2021;USA
Chevrolet;Malibu;27.0;6;2500;240;2900;2022;USA
Toyota;Camry;34.0;4;2500;200;2900;2023;Japan
Honda;Civic;35.0;4;1800;140;2600;2022;Japan
BMW;X5;24.0;8;4000;450;4000;2023;Germany
Mercedes-Benz;E-Class;28.0;6;3000;340;3200;2022;Germany
Hyundai;Sonata;32.0;4;2400;190;2800;2023;South Korea
Nissan;Maxima;28.5;6;3000;290;3100;2022;Japan
Audi;Q5;26.0;6;3200;350;3300;2022;Germany
Lexus;RX;31.0;6;3500;300;3400;2023;Japan
Kia;Sorento;25.0;4;2400;200;3000;2022;South Korea
Subaru;Outback;33.5;6;3300;260;3100;2023;Japan
Volkswagen;Jetta;30.5;4;2600;220;2800;2022;Germany
Mazda;CX-5;29.0;4;2500;210;2900;2022;Japan
Tesla;Model S;120.0;0;0;500;3800;2023;USA